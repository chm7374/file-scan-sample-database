This is an executable file of a programming language!
